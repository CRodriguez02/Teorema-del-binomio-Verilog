module SUM(
input  [31:0] op1, op2,
output [31:0] SUMA 
);


assign SUMA=op1+op2;

endmodule 