module SUM_4(
input  [31:0] op1,
output [31:0] SUMA 
);


assign SUMA=op1+9'd4;

endmodule 