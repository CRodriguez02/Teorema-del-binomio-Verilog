module mult5(
input in_and,
input [31:0] in_x, in_y,
output reg [31:0] out_z
);
always@(*)
begin 
	case (in_and)
		1'b0:
			begin
				out_z=in_x;
			end
		1'b1:
			begin
				out_z=in_y;
			end
		endcase
	end

endmodule 