module MA(
input  op1,op2,
output AND
);

assign AND=op1&op2;

endmodule 